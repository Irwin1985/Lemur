module ast

pub interface Node {
	to_string() string
}