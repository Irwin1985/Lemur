module ast

pub struct None {
	
}

fn (n None) to_string() string {
	return ""
}